SRAM (single-port)

ONE array

ONE port → read OR write
-----------------------------------------------------------
-----------------------------------------------------------
Simple DPRAM

ONE array

Port A = write

Port B = read
-----------------------------------------------------------
-----------------------------------------------------------
True DPRAM

ONE array

Port A = read/write

Port B = read/write
